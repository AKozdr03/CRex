/**
 * KK & AK Company
 * 
 * Authors: Krzysztof Korbaś, Andrzej Kozdrowski
 * 
 * Description:
 * Top console module.
 **/

module top_console(


    );
    
    
endmodule