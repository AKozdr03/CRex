/**
 * KK & AK Company
 * 
 * Authors: Krzysztof Korbaś, Andrzej Kozdrowski
 * 
 * Description:
 * Testbench of top console module.
 **/

module top_console_tb();
    
    
    
endmodule