/**
 * KK & AK Company
 * 
 * Authors: Krzysztof Korbaś, Andrzej Kozdrowski
 * 
 * Description:
 * Top fpga module.
 **/

module top_fpga(


);



endmodule